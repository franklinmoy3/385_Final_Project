
module spriteTable(input logic clk,
							output logic [0:24][0:17][0:5] blueTank,
							output logic [0:24][0:17][0:5] redTank,
							);

always_comb
begin

blueTank <=
'{
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,0,1,1,5,0,0,0,0,0,0,0},
'{0,0,0,0,11,0,0,0,3,3,0,0,0,11,0,0,0,0},
'{0,0,8,15,10,14,14,15,2,1,15,14,14,14,11,8,8,0},
'{0,8,5,8,15,14,14,15,2,1,15,14,14,15,8,5,8,0},
'{0,8,8,8,0,11,15,15,2,1,15,15,11,0,8,8,8,0},
'{0,8,5,5,8,15,14,11,2,1,11,14,15,8,5,5,5,0},
'{0,8,5,5,8,14,14,11,2,1,11,14,14,8,8,5,8,0},
'{0,8,5,8,11,10,14,11,2,1,11,14,14,11,8,8,8,0},
'{0,8,5,8,14,14,10,15,3,2,11,10,14,14,8,5,8,0},
'{0,8,8,8,14,10,14,11,9,9,11,14,10,14,15,8,8,0},
'{0,8,8,15,14,14,14,10,12,10,14,14,14,14,15,8,8,0},
'{0,0,15,11,14,14,14,14,10,10,14,14,14,14,11,15,0,0},
'{0,8,11,11,14,14,11,3,2,2,3,11,14,14,11,11,8,0},
'{0,0,11,11,14,14,11,11,14,14,11,11,14,14,11,11,0,0},
'{0,8,11,14,14,14,14,11,11,11,11,14,14,14,11,14,8,0},
'{0,0,14,14,15,14,14,11,2,11,14,14,14,13,14,14,0,0},
'{0,0,11,14,15,11,14,11,4,11,14,14,11,15,14,14,8,0},
'{0,0,11,14,15,15,11,11,11,14,14,11,15,15,11,14,0,0},
'{0,0,11,14,15,15,2,3,15,15,3,2,15,15,14,14,8,0},
'{0,8,11,14,15,13,11,11,11,11,11,15,13,15,14,11,8,0},
'{0,0,8,11,14,13,0,0,11,11,0,0,15,14,11,8,0,0},
'{0,0,0,13,11,0,0,0,0,0,0,0,15,13,11,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};

red <=
'{
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,4,1,1,0,0,0,0,0,0,0,0},
'{0,0,0,0,0,0,0,4,1,2,0,0,0,0,0,0,0,0},
'{0,0,0,0,15,0,0,0,2,3,0,0,11,15,0,0,0,0},
'{0,8,0,15,9,9,15,12,1,2,12,14,9,9,11,8,0,0},
'{0,8,5,8,11,10,15,11,1,2,11,14,9,11,8,5,8,0},
'{0,8,8,8,0,15,11,11,1,2,12,11,15,0,8,8,8,0},
'{0,5,5,5,0,11,14,11,1,2,15,14,11,8,5,5,8,0},
'{0,8,5,8,0,10,14,11,1,2,11,9,14,0,5,5,8,0},
'{0,8,8,0,15,9,14,11,1,2,11,14,9,11,8,5,8,0},
'{0,8,5,8,14,10,14,12,2,3,12,14,10,14,8,5,8,0},
'{0,8,8,11,14,9,15,15,9,9,15,14,10,14,8,8,8,0},
'{0,8,8,11,14,10,15,9,9,9,14,15,10,14,12,8,8,0},
'{0,8,11,15,14,14,15,9,9,9,14,15,14,14,15,11,0,0},
'{0,8,15,15,14,15,11,6,6,6,6,11,14,14,15,15,8,0},
'{0,0,15,15,14,14,11,15,15,15,15,11,14,14,15,11,0,0},
'{0,8,14,15,15,14,15,15,15,15,11,14,14,15,15,15,8,0},
'{0,0,14,14,11,15,14,6,3,15,14,14,15,11,14,15,0,0},
'{0,8,14,14,11,15,15,11,8,15,13,15,11,11,14,15,0,0},
'{0,0,15,15,11,11,15,15,15,14,15,5,11,11,15,15,0,0},
'{0,0,14,14,11,8,2,6,11,11,3,3,11,11,14,15,0,0},
'{0,8,15,14,11,11,11,15,15,15,15,11,11,11,10,15,8,0},
'{0,0,12,15,14,11,0,0,0,0,0,0,15,14,15,0,0,0},
'{0,0,0,15,15,0,0,0,0,0,0,0,12,15,15,0,0,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
};

end

endmodule